library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package dat_t_pkg is

	type dat_t is array(7 downto 0) of std_logic_vector;
	
end package dat_t_pkg;