library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity back_fsm is
	port (
		bvalid	:	out std_logic;		-- data valid / ready to load
		bload		:	in std_logic;		-- load data / send acknowledge
		b_en		:	in std_logic;		-- enable receipt of adata
		bclk		:	in std_logic;
		brst_n	:	in std_logic
	);
end entity back_fsm;

architecture RTL of back_fsm is
	type state_t is (READY, ESPERA);
	signal state, next_state : state_t;
begin
	-- State register
	process (bclk, brst_n)
	begin
		if (brst_n = '0') then
			state <= ESPERA;
		elsif (rising_edge(bclk)) then
			state <= next_state;
		end if;
	end process;

	-- Next state logic
	process (state, bload, b_en)
	begin
		case state is
			when READY =>
				if (bload = '1') then
					next_state <= ESPERA;
				else
					next_state <= READY;
				end if;
			when ESPERA =>
				if (b_en = '1') then
					next_state <= READY;
				else
					next_state <= ESPERA;
				end if;
		end case;
	end process;

	-- Output assignment
	bvalid <= '1' when state = READY else '0';
end architecture RTL;